magic
tech sky130A
timestamp 1689005540
<< nwell >>
rect -950 200 1900 1100
rect -950 -1950 1900 -1100
<< nmos >>
rect -500 -250 -450 -50
rect 200 -250 250 -50
rect 900 -250 950 -50
rect 1600 -250 1650 -50
rect -500 -750 -450 -550
rect 200 -750 250 -550
rect 900 -750 950 -550
rect -500 -2400 -450 -2200
rect 0 -2400 50 -2200
rect 900 -2400 950 -2200
rect 1600 -2400 1650 -2200
rect -500 -2850 -450 -2650
<< pmos >>
rect -500 650 -450 850
rect -500 250 -450 450
rect 200 250 250 450
rect 900 250 950 450
rect 1600 250 1650 450
rect -500 -1400 -450 -1200
rect -500 -1900 -450 -1700
rect 0 -1900 50 -1700
rect 900 -1900 950 -1700
rect 1600 -1900 1650 -1700
<< ndiff >>
rect -700 -100 -500 -50
rect -700 -200 -650 -100
rect -550 -200 -500 -100
rect -700 -250 -500 -200
rect -450 -100 -250 -50
rect -450 -200 -400 -100
rect -300 -200 -250 -100
rect -450 -250 -250 -200
rect 0 -100 200 -50
rect 0 -200 50 -100
rect 150 -200 200 -100
rect 0 -250 200 -200
rect 250 -100 450 -50
rect 250 -200 300 -100
rect 400 -200 450 -100
rect 250 -250 450 -200
rect 700 -100 900 -50
rect 700 -200 750 -100
rect 850 -200 900 -100
rect 700 -250 900 -200
rect 950 -100 1150 -50
rect 950 -200 1000 -100
rect 1100 -200 1150 -100
rect 950 -250 1150 -200
rect 1400 -100 1600 -50
rect 1400 -200 1450 -100
rect 1550 -200 1600 -100
rect 1400 -250 1600 -200
rect 1650 -100 1850 -50
rect 1650 -200 1700 -100
rect 1800 -200 1850 -100
rect 1650 -250 1850 -200
rect -700 -600 -500 -550
rect -700 -700 -650 -600
rect -550 -700 -500 -600
rect -700 -750 -500 -700
rect -450 -600 -250 -550
rect -450 -700 -400 -600
rect -300 -700 -250 -600
rect -450 -750 -250 -700
rect 0 -600 200 -550
rect 0 -700 50 -600
rect 150 -700 200 -600
rect 0 -750 200 -700
rect 250 -600 450 -550
rect 250 -700 300 -600
rect 400 -700 450 -600
rect 250 -750 450 -700
rect 700 -600 900 -550
rect 700 -700 750 -600
rect 850 -700 900 -600
rect 700 -750 900 -700
rect 950 -600 1150 -550
rect 950 -700 1000 -600
rect 1100 -700 1150 -600
rect 950 -750 1150 -700
rect -700 -2250 -500 -2200
rect -700 -2350 -650 -2250
rect -550 -2350 -500 -2250
rect -700 -2400 -500 -2350
rect -450 -2250 -250 -2200
rect -450 -2350 -400 -2250
rect -300 -2350 -250 -2250
rect -450 -2400 -250 -2350
rect -200 -2250 0 -2200
rect -200 -2350 -150 -2250
rect -50 -2350 0 -2250
rect -200 -2400 0 -2350
rect 50 -2250 250 -2200
rect 50 -2350 100 -2250
rect 200 -2350 250 -2250
rect 50 -2400 250 -2350
rect 700 -2250 900 -2200
rect 700 -2350 750 -2250
rect 850 -2350 900 -2250
rect 700 -2400 900 -2350
rect 950 -2250 1150 -2200
rect 950 -2350 1000 -2250
rect 1100 -2350 1150 -2250
rect 950 -2400 1150 -2350
rect 1400 -2250 1600 -2200
rect 1400 -2350 1450 -2250
rect 1550 -2350 1600 -2250
rect 1400 -2400 1600 -2350
rect 1650 -2250 1850 -2200
rect 1650 -2350 1700 -2250
rect 1800 -2350 1850 -2250
rect 1650 -2400 1850 -2350
rect -700 -2700 -500 -2650
rect -700 -2800 -650 -2700
rect -550 -2800 -500 -2700
rect -700 -2850 -500 -2800
rect -450 -2700 -250 -2650
rect -450 -2800 -400 -2700
rect -300 -2800 -250 -2700
rect -450 -2850 -250 -2800
<< pdiff >>
rect -700 800 -500 850
rect -700 700 -650 800
rect -550 700 -500 800
rect -700 650 -500 700
rect -450 800 -250 850
rect -450 700 -400 800
rect -300 700 -250 800
rect -450 650 -250 700
rect -700 400 -500 450
rect -700 300 -650 400
rect -550 300 -500 400
rect -700 250 -500 300
rect -450 400 -250 450
rect -450 300 -400 400
rect -300 300 -250 400
rect -450 250 -250 300
rect 0 400 200 450
rect 0 300 50 400
rect 150 300 200 400
rect 0 250 200 300
rect 250 400 450 450
rect 250 300 300 400
rect 400 300 450 400
rect 250 250 450 300
rect 700 400 900 450
rect 700 300 750 400
rect 850 300 900 400
rect 700 250 900 300
rect 950 400 1150 450
rect 950 300 1000 400
rect 1100 300 1150 400
rect 950 250 1150 300
rect 1400 400 1600 450
rect 1400 300 1450 400
rect 1550 300 1600 400
rect 1400 250 1600 300
rect 1650 400 1850 450
rect 1650 300 1700 400
rect 1800 300 1850 400
rect 1650 250 1850 300
rect -700 -1250 -500 -1200
rect -700 -1350 -650 -1250
rect -550 -1350 -500 -1250
rect -700 -1400 -500 -1350
rect -450 -1250 -250 -1200
rect -450 -1350 -400 -1250
rect -300 -1350 -250 -1250
rect -450 -1400 -250 -1350
rect -700 -1750 -500 -1700
rect -700 -1850 -650 -1750
rect -550 -1850 -500 -1750
rect -700 -1900 -500 -1850
rect -450 -1750 -250 -1700
rect -450 -1850 -400 -1750
rect -300 -1850 -250 -1750
rect -450 -1900 -250 -1850
rect -200 -1750 0 -1700
rect -200 -1850 -150 -1750
rect -50 -1850 0 -1750
rect -200 -1900 0 -1850
rect 50 -1750 250 -1700
rect 50 -1850 100 -1750
rect 200 -1850 250 -1750
rect 50 -1900 250 -1850
rect 700 -1750 900 -1700
rect 700 -1850 750 -1750
rect 850 -1850 900 -1750
rect 700 -1900 900 -1850
rect 950 -1750 1150 -1700
rect 950 -1850 1000 -1750
rect 1100 -1850 1150 -1750
rect 950 -1900 1150 -1850
rect 1400 -1750 1600 -1700
rect 1400 -1850 1450 -1750
rect 1550 -1850 1600 -1750
rect 1400 -1900 1600 -1850
rect 1650 -1750 1850 -1700
rect 1650 -1850 1700 -1750
rect 1800 -1850 1850 -1750
rect 1650 -1900 1850 -1850
<< ndiffc >>
rect -650 -200 -550 -100
rect -400 -200 -300 -100
rect 50 -200 150 -100
rect 300 -200 400 -100
rect 750 -200 850 -100
rect 1000 -200 1100 -100
rect 1450 -200 1550 -100
rect 1700 -200 1800 -100
rect -650 -700 -550 -600
rect -400 -700 -300 -600
rect 50 -700 150 -600
rect 300 -700 400 -600
rect 750 -700 850 -600
rect 1000 -700 1100 -600
rect -650 -2350 -550 -2250
rect -400 -2350 -300 -2250
rect -150 -2350 -50 -2250
rect 100 -2350 200 -2250
rect 750 -2350 850 -2250
rect 1000 -2350 1100 -2250
rect 1450 -2350 1550 -2250
rect 1700 -2350 1800 -2250
rect -650 -2800 -550 -2700
rect -400 -2800 -300 -2700
<< pdiffc >>
rect -650 700 -550 800
rect -400 700 -300 800
rect -650 300 -550 400
rect -400 300 -300 400
rect 50 300 150 400
rect 300 300 400 400
rect 750 300 850 400
rect 1000 300 1100 400
rect 1450 300 1550 400
rect 1700 300 1800 400
rect -650 -1350 -550 -1250
rect -400 -1350 -300 -1250
rect -650 -1850 -550 -1750
rect -400 -1850 -300 -1750
rect -150 -1850 -50 -1750
rect 100 -1850 200 -1750
rect 750 -1850 850 -1750
rect 1000 -1850 1100 -1750
rect 1450 -1850 1550 -1750
rect 1700 -1850 1800 -1750
<< psubdiff >>
rect -900 -100 -700 -50
rect -900 -200 -850 -100
rect -750 -200 -700 -100
rect -900 -250 -700 -200
rect -200 -100 0 -50
rect -200 -200 -150 -100
rect -50 -200 0 -100
rect -200 -250 0 -200
rect 500 -100 700 -50
rect 500 -200 550 -100
rect 650 -200 700 -100
rect 500 -250 700 -200
rect 1200 -150 1400 -50
rect 1200 -200 1250 -150
rect 1300 -200 1400 -150
rect 1200 -250 1400 -200
rect -900 -600 -700 -550
rect -900 -700 -850 -600
rect -750 -700 -700 -600
rect -900 -750 -700 -700
rect -200 -600 0 -550
rect -200 -700 -150 -600
rect -50 -700 0 -600
rect -200 -750 0 -700
rect 500 -600 700 -550
rect 500 -700 550 -600
rect 650 -700 700 -600
rect 500 -750 700 -700
rect -900 -2250 -700 -2200
rect -900 -2350 -850 -2250
rect -750 -2350 -700 -2250
rect -900 -2400 -700 -2350
rect 500 -2250 700 -2200
rect 500 -2350 550 -2250
rect 650 -2350 700 -2250
rect 500 -2400 700 -2350
rect 1200 -2250 1400 -2200
rect 1200 -2350 1250 -2250
rect 1350 -2350 1400 -2250
rect 1200 -2400 1400 -2350
rect -900 -2700 -700 -2650
rect -900 -2800 -850 -2700
rect -750 -2800 -700 -2700
rect -900 -2850 -700 -2800
<< nsubdiff >>
rect -900 800 -700 850
rect -900 700 -850 800
rect -750 700 -700 800
rect -900 650 -700 700
rect -900 400 -700 450
rect -900 300 -850 400
rect -750 300 -700 400
rect -900 250 -700 300
rect -200 400 0 450
rect -200 300 -150 400
rect -50 300 0 400
rect -200 250 0 300
rect 500 400 700 450
rect 500 300 550 400
rect 650 300 700 400
rect 500 250 700 300
rect 1200 400 1400 450
rect 1200 300 1250 400
rect 1350 300 1400 400
rect 1200 250 1400 300
rect -900 -1250 -700 -1200
rect -900 -1350 -850 -1250
rect -750 -1350 -700 -1250
rect -900 -1400 -700 -1350
rect 500 -1750 700 -1700
rect 500 -1850 550 -1750
rect 650 -1850 700 -1750
rect 500 -1900 700 -1850
rect 1200 -1750 1400 -1700
rect 1200 -1850 1250 -1750
rect 1350 -1850 1400 -1750
rect 1200 -1900 1400 -1850
<< psubdiffcont >>
rect -850 -200 -750 -100
rect -150 -200 -50 -100
rect 550 -200 650 -100
rect 1250 -200 1300 -150
rect -850 -700 -750 -600
rect -150 -700 -50 -600
rect 550 -700 650 -600
rect -850 -2350 -750 -2250
rect 550 -2350 650 -2250
rect 1250 -2350 1350 -2250
rect -850 -2800 -750 -2700
<< nsubdiffcont >>
rect -850 700 -750 800
rect -850 300 -750 400
rect -150 300 -50 400
rect 550 300 650 400
rect 1250 300 1350 400
rect -850 -1350 -750 -1250
rect 550 -1850 650 -1750
rect 1250 -1850 1350 -1750
<< poly >>
rect -500 1000 -350 1050
rect -500 950 -450 1000
rect -400 950 -350 1000
rect -500 900 -350 950
rect -500 850 -450 900
rect -500 600 -450 650
rect 900 600 1050 650
rect 900 550 950 600
rect 1000 550 1050 600
rect 900 500 1050 550
rect 1600 600 1750 650
rect 1600 550 1650 600
rect 1700 550 1750 600
rect 1600 500 1750 550
rect -500 450 -450 500
rect 200 450 250 500
rect 900 450 950 500
rect 1600 450 1650 500
rect -750 100 -600 150
rect -500 100 -450 250
rect -750 50 -700 100
rect -650 50 -450 100
rect -750 0 -600 50
rect -500 -50 -450 50
rect 200 -50 250 250
rect 900 200 950 250
rect 1600 200 1650 250
rect 800 100 950 150
rect 800 50 850 100
rect 900 50 950 100
rect 800 0 950 50
rect 1550 100 1700 150
rect 1550 50 1600 100
rect 1650 50 1700 100
rect 1550 0 1700 50
rect 900 -50 950 0
rect 1600 -50 1650 0
rect -500 -300 -450 -250
rect 200 -300 250 -250
rect 900 -300 950 -250
rect 1600 -300 1650 -250
rect 100 -350 250 -300
rect 100 -400 150 -350
rect 200 -400 250 -350
rect 100 -450 250 -400
rect -500 -550 -450 -500
rect 200 -550 250 -500
rect 900 -550 950 -500
rect 1250 -600 1400 -550
rect 1250 -650 1300 -600
rect 1350 -650 1400 -600
rect 1250 -700 1400 -650
rect -500 -800 -450 -750
rect 200 -800 250 -750
rect -600 -850 -450 -800
rect -900 -900 -750 -850
rect -900 -950 -850 -900
rect -800 -950 -750 -900
rect -600 -900 -550 -850
rect -500 -900 -450 -850
rect -600 -950 -450 -900
rect 100 -850 250 -800
rect 900 -800 950 -750
rect 1250 -800 1300 -700
rect 900 -850 1350 -800
rect 100 -900 150 -850
rect 200 -900 250 -850
rect 100 -950 250 -900
rect 1200 -900 1250 -850
rect 1300 -900 1350 -850
rect 1200 -950 1350 -900
rect -900 -1000 -750 -950
rect -850 -1100 -800 -1000
rect -850 -1150 -450 -1100
rect -500 -1200 -450 -1150
rect -500 -1450 -450 -1400
rect -500 -1700 -450 -1650
rect 0 -1700 50 -1650
rect 900 -1700 950 -1650
rect 1600 -1700 1650 -1650
rect -700 -2050 -550 -2000
rect -500 -2050 -450 -1900
rect -700 -2100 -650 -2050
rect -600 -2100 -450 -2050
rect -700 -2150 -550 -2100
rect -500 -2200 -450 -2100
rect -200 -2050 -50 -2000
rect 0 -2050 50 -1900
rect -200 -2100 -150 -2050
rect -100 -2100 50 -2050
rect -200 -2150 -50 -2100
rect 0 -2200 50 -2100
rect 700 -2050 850 -2000
rect 900 -2050 950 -1900
rect 700 -2100 750 -2050
rect 800 -2100 950 -2050
rect 700 -2150 850 -2100
rect 900 -2200 950 -2100
rect 1350 -2050 1500 -2000
rect 1600 -2050 1650 -1900
rect 1350 -2100 1400 -2050
rect 1450 -2100 1650 -2050
rect 1350 -2150 1500 -2100
rect 1600 -2200 1650 -2100
rect -500 -2450 -450 -2400
rect 0 -2450 50 -2400
rect 900 -2450 950 -2400
rect 1600 -2450 1650 -2400
rect -500 -2650 -450 -2600
rect -500 -2900 -450 -2850
rect -900 -2950 -450 -2900
rect -900 -3000 -850 -2950
rect -800 -3000 -750 -2950
rect -900 -3050 -750 -3000
<< polycont >>
rect -450 950 -400 1000
rect 950 550 1000 600
rect 1650 550 1700 600
rect -700 50 -650 100
rect 850 50 900 100
rect 1600 50 1650 100
rect 150 -400 200 -350
rect 1300 -650 1350 -600
rect -850 -950 -800 -900
rect -550 -900 -500 -850
rect 150 -900 200 -850
rect 1250 -900 1300 -850
rect -650 -2100 -600 -2050
rect -150 -2100 -100 -2050
rect 750 -2100 800 -2050
rect 1400 -2100 1450 -2050
rect -850 -3000 -800 -2950
<< locali >>
rect -18000 12000 -8000 13000
rect -18000 4000 -17000 12000
rect -9000 4000 -8000 12000
rect -18000 3000 -8000 4000
rect -5000 12000 5000 13000
rect -5000 4000 -4000 12000
rect 4000 4000 5000 12000
rect -5000 3000 5000 4000
rect 8000 12000 18000 13000
rect 8000 4000 9000 12000
rect 17000 4000 18000 12000
rect 8000 3000 18000 4000
rect 12650 2450 14050 2500
rect 750 1500 1000 1550
rect 750 1350 800 1500
rect 950 1350 1000 1500
rect 750 1300 1000 1350
rect 12650 1250 12700 2450
rect 14000 1250 14050 2450
rect 12650 1200 14050 1250
rect -500 1000 -350 1050
rect -500 950 -450 1000
rect -400 950 -350 1000
rect -500 900 -350 950
rect -900 800 -700 850
rect 500 800 700 850
rect -900 700 -850 800
rect -750 700 -650 800
rect -550 700 -500 800
rect -450 700 -400 800
rect -300 700 150 800
rect -900 650 -700 700
rect -850 400 -750 650
rect -150 600 0 650
rect -150 550 -100 600
rect -50 550 0 600
rect -150 500 0 550
rect -850 250 -750 300
rect -700 400 -500 450
rect -150 400 -50 500
rect 50 450 150 700
rect 500 700 550 800
rect 650 700 700 800
rect 500 650 700 700
rect 1250 650 1400 700
rect 550 450 650 650
rect 900 600 1300 650
rect 1350 600 1750 650
rect 900 550 950 600
rect 1000 550 1650 600
rect 1700 550 1750 600
rect 900 500 1050 550
rect 1600 500 1750 550
rect -700 300 -650 400
rect -550 300 -500 400
rect -450 300 -400 400
rect -300 300 -250 400
rect -700 250 -500 300
rect -750 100 -600 150
rect -750 50 -700 100
rect -650 50 -600 100
rect -750 0 -600 50
rect -400 -50 -300 300
rect -150 250 -50 300
rect 0 400 200 450
rect 500 400 700 450
rect 1200 400 1400 450
rect 0 300 50 400
rect 150 300 200 400
rect 250 300 300 400
rect 400 300 450 400
rect 500 300 550 400
rect 650 300 750 400
rect 850 300 900 400
rect 950 300 1000 400
rect 1100 300 1150 400
rect 1200 300 1250 400
rect 1350 300 1450 400
rect 1550 300 1600 400
rect 1650 300 1700 400
rect 1800 300 1850 400
rect 0 250 200 300
rect 300 150 400 300
rect 500 250 700 300
rect 300 100 450 150
rect 300 50 350 100
rect 400 50 450 100
rect 300 0 450 50
rect 800 100 950 150
rect 800 50 850 100
rect 900 50 950 100
rect 800 0 950 50
rect -450 -100 -250 -50
rect 300 -100 400 0
rect 1000 -50 1100 300
rect 1200 250 1400 300
rect 1550 100 1700 150
rect 1550 50 1600 100
rect 1650 50 1700 100
rect 1550 0 1700 50
rect 1750 -50 1850 300
rect 500 -100 700 -50
rect -900 -200 -850 -100
rect -750 -200 -650 -100
rect -550 -200 -500 -100
rect -450 -200 -400 -100
rect -300 -200 -250 -100
rect -200 -200 -150 -100
rect -50 -200 50 -100
rect 150 -200 200 -100
rect 250 -200 300 -100
rect 400 -200 450 -100
rect 500 -200 550 -100
rect 650 -200 700 -100
rect -450 -250 -250 -200
rect -400 -300 -300 -250
rect -400 -350 250 -300
rect -400 -400 150 -350
rect 200 -400 250 -350
rect 100 -450 250 -400
rect -1000 -600 -700 -550
rect -450 -600 -250 -550
rect 300 -600 400 -200
rect 500 -250 700 -200
rect 750 -100 850 -50
rect 750 -350 850 -200
rect 950 -100 1150 -50
rect 950 -200 1000 -100
rect 1100 -200 1150 -100
rect 950 -250 1150 -200
rect 1200 -150 1400 -50
rect 1200 -200 1250 -150
rect 1300 -200 1400 -150
rect 1200 -250 1400 -200
rect 1450 -100 1550 -50
rect 1450 -350 1550 -200
rect 1650 -100 1850 -50
rect 1650 -200 1700 -100
rect 1800 -200 1850 -100
rect 1650 -250 1850 -200
rect 750 -450 1550 -350
rect 500 -600 700 -550
rect 1000 -600 1100 -450
rect 1250 -600 1400 -550
rect -1000 -650 -850 -600
rect -900 -700 -850 -650
rect -750 -700 -650 -600
rect -550 -700 -500 -600
rect -450 -700 -400 -600
rect -300 -700 -250 -600
rect -200 -700 -150 -600
rect -50 -700 50 -600
rect 150 -700 200 -600
rect 250 -700 300 -600
rect 400 -700 450 -600
rect 500 -700 550 -600
rect 650 -700 750 -600
rect 850 -700 900 -600
rect 950 -700 1000 -600
rect 1100 -700 1150 -600
rect 1250 -650 1300 -600
rect 1350 -650 1400 -600
rect 1250 -700 1400 -650
rect 1450 -700 1600 -650
rect -900 -750 -700 -700
rect -450 -750 -250 -700
rect 300 -750 400 -700
rect 500 -750 700 -700
rect 1000 -750 1100 -700
rect 1450 -750 1500 -700
rect 1550 -750 1600 -700
rect -600 -850 -450 -800
rect -900 -900 -750 -850
rect -900 -950 -850 -900
rect -800 -950 -750 -900
rect -600 -900 -550 -850
rect -500 -900 -450 -850
rect -600 -950 -450 -900
rect -900 -1000 -750 -950
rect -400 -1000 -300 -750
rect 1450 -800 1600 -750
rect 1700 -800 1800 -250
rect 2050 -650 2100 -550
rect 100 -850 250 -800
rect 100 -900 150 -850
rect 200 -900 250 -850
rect 100 -950 250 -900
rect 1200 -850 1350 -800
rect 1200 -900 1250 -850
rect 1300 -900 1350 -850
rect 1200 -950 1350 -900
rect 1650 -850 1800 -800
rect 1650 -900 1700 -850
rect 1750 -900 1800 -850
rect 1650 -950 1800 -900
rect -400 -1100 400 -1000
rect -700 -1250 -500 -1200
rect -900 -1350 -850 -1250
rect -750 -1350 -650 -1250
rect -550 -1350 -500 -1250
rect -700 -1400 -500 -1350
rect -400 -1250 -300 -1200
rect -400 -1500 -300 -1350
rect 300 -1450 400 -1100
rect 700 -1250 900 -1200
rect 700 -1350 750 -1250
rect 850 -1350 900 -1250
rect 700 -1400 900 -1350
rect 1250 -1300 1350 -950
rect 1250 -1350 1800 -1300
rect 1250 -1400 1700 -1350
rect 1750 -1400 1800 -1350
rect 250 -1500 450 -1450
rect -650 -1600 -50 -1500
rect -650 -1700 -550 -1600
rect -150 -1700 -50 -1600
rect 250 -1600 300 -1500
rect 400 -1600 450 -1500
rect 250 -1650 450 -1600
rect -700 -1750 -500 -1700
rect -700 -1850 -650 -1750
rect -550 -1850 -500 -1750
rect -700 -1900 -500 -1850
rect -400 -1750 -300 -1700
rect -400 -2000 -300 -1850
rect -200 -1750 0 -1700
rect -200 -1850 -150 -1750
rect -50 -1850 0 -1750
rect -200 -1900 0 -1850
rect 100 -1750 200 -1700
rect 750 -1750 850 -1400
rect 1650 -1450 1800 -1400
rect 1250 -1600 1950 -1500
rect 1250 -1750 1350 -1600
rect 1850 -1650 1950 -1600
rect 1450 -1750 1550 -1700
rect 500 -1850 550 -1750
rect 650 -1850 750 -1750
rect 850 -1850 900 -1750
rect 950 -1850 1000 -1750
rect 1100 -1850 1150 -1750
rect 1350 -1850 1450 -1750
rect -700 -2050 -550 -2000
rect -700 -2100 -650 -2050
rect -600 -2100 -550 -2050
rect -700 -2150 -550 -2100
rect -400 -2050 -250 -2000
rect -400 -2100 -350 -2050
rect -300 -2100 -250 -2050
rect -400 -2150 -250 -2100
rect -200 -2050 -50 -2000
rect -200 -2100 -150 -2050
rect -100 -2100 -50 -2050
rect -200 -2150 -50 -2100
rect -1000 -2250 -750 -2150
rect -400 -2250 -300 -2150
rect 100 -2200 200 -1850
rect 700 -2050 850 -2000
rect 700 -2100 750 -2050
rect 800 -2100 850 -2050
rect 700 -2150 850 -2100
rect -150 -2250 -50 -2200
rect 50 -2250 250 -2200
rect 1000 -2250 1100 -1850
rect 1250 -1900 1350 -1850
rect 1450 -1900 1550 -1850
rect 1700 -1750 1800 -1700
rect 1350 -2050 1500 -2000
rect 1350 -2100 1400 -2050
rect 1450 -2100 1500 -2050
rect 1350 -2150 1500 -2100
rect 1700 -2250 1800 -1850
rect -700 -2350 -650 -2250
rect -550 -2350 -500 -2250
rect -450 -2350 -400 -2250
rect -300 -2350 -250 -2250
rect -200 -2350 -150 -2250
rect -50 -2350 0 -2250
rect 50 -2350 100 -2250
rect 200 -2350 250 -2250
rect 450 -2350 550 -2250
rect 650 -2350 750 -2250
rect 850 -2350 900 -2250
rect 950 -2350 1000 -2250
rect 1100 -2350 1150 -2250
rect 1200 -2350 1250 -2250
rect 1350 -2350 1450 -2250
rect 1550 -2350 1600 -2250
rect -850 -2400 -750 -2350
rect -650 -2450 -550 -2350
rect -150 -2450 -50 -2350
rect 50 -2400 250 -2350
rect -650 -2550 -50 -2450
rect -1000 -2650 -750 -2550
rect -850 -2700 -750 -2650
rect -650 -2700 -550 -2650
rect -900 -2800 -850 -2700
rect -750 -2800 -650 -2700
rect -650 -2850 -550 -2800
rect -400 -2700 -300 -2550
rect -400 -2850 -300 -2800
rect -900 -2950 -750 -2900
rect -900 -3000 -850 -2950
rect -800 -3000 -750 -2950
rect -1000 -3050 -950 -3000
rect -900 -3050 -750 -3000
rect -1100 -3100 -950 -3050
rect 550 -3100 650 -2350
rect 1000 -2800 1100 -2350
rect 950 -2850 1150 -2800
rect 950 -2950 1000 -2850
rect 1100 -2950 1150 -2850
rect 950 -3000 1150 -2950
rect 1400 -3100 1500 -2350
rect 1700 -2400 1800 -2350
rect -1100 -3150 1500 -3100
rect -1000 -3200 1500 -3150
rect -18000 -6000 -8000 -5000
rect -18000 -14000 -17000 -6000
rect -9000 -14000 -8000 -6000
rect -18000 -15000 -8000 -14000
rect -5000 -6000 5000 -5000
rect -5000 -14000 -4000 -6000
rect 4000 -14000 5000 -6000
rect -5000 -15000 5000 -14000
rect 8000 -6000 18000 -5000
rect 8000 -14000 9000 -6000
rect 17000 -14000 18000 -6000
rect 8000 -15000 18000 -14000
<< viali >>
rect -17000 4000 -9000 12000
rect -4000 4000 4000 12000
rect 9000 4000 17000 12000
rect 800 1350 950 1500
rect 12700 1250 14000 2450
rect -1100 950 -1000 1050
rect -450 950 -400 1000
rect 1950 950 2050 1050
rect -1100 750 -1000 850
rect -850 700 -750 800
rect -1100 550 -1000 650
rect -1100 350 -1000 450
rect -100 550 -50 600
rect 550 700 650 800
rect 1950 750 2050 850
rect 1300 600 1350 650
rect 1950 550 2050 650
rect -650 300 -550 400
rect -1100 150 -1000 250
rect -700 50 -650 100
rect -1100 -50 -1000 50
rect 50 300 150 400
rect 550 300 650 400
rect 1250 300 1350 400
rect 1950 350 2050 450
rect 350 50 400 100
rect 850 50 900 100
rect 1600 50 1650 100
rect 1950 150 2050 250
rect 1950 -50 2050 50
rect -1100 -250 -1000 -150
rect -850 -200 -750 -100
rect -400 -200 -300 -100
rect 50 -200 150 -100
rect 550 -200 650 -100
rect -1100 -450 -1000 -350
rect -1100 -650 -1000 -550
rect 1000 -200 1100 -100
rect 1250 -200 1300 -150
rect 1700 -200 1800 -100
rect 1950 -250 2050 -150
rect -850 -700 -750 -600
rect -400 -700 -300 -600
rect 50 -700 150 -600
rect 550 -700 650 -600
rect 1300 -650 1350 -600
rect 1500 -750 1550 -700
rect -1100 -850 -1000 -750
rect -850 -950 -800 -900
rect -550 -900 -500 -850
rect -1100 -1050 -1000 -950
rect 1950 -450 2050 -350
rect 1950 -650 2050 -550
rect 150 -900 200 -850
rect 1950 -850 2050 -750
rect 1700 -900 1750 -850
rect -1100 -1250 -1000 -1150
rect -650 -1350 -550 -1250
rect -1100 -1450 -1000 -1350
rect 750 -1350 850 -1250
rect 1950 -1050 2050 -950
rect 1950 -1250 2050 -1150
rect 1700 -1400 1750 -1350
rect -1100 -1650 -1000 -1550
rect 300 -1600 400 -1500
rect -1100 -1850 -1000 -1750
rect -1100 -2050 -1000 -1950
rect 1950 -1450 2050 -1350
rect 1950 -1650 2050 -1550
rect -650 -2100 -600 -2050
rect -350 -2100 -300 -2050
rect -150 -2100 -100 -2050
rect -1100 -2250 -1000 -2150
rect 750 -2100 800 -2050
rect 1700 -1850 1800 -1750
rect 1950 -1850 2050 -1750
rect 1400 -2100 1450 -2050
rect 1950 -2050 2050 -1950
rect 1950 -2250 2050 -2150
rect 100 -2350 200 -2250
rect -1100 -2450 -1000 -2350
rect -1100 -2650 -1000 -2550
rect -1100 -2850 -1000 -2750
rect -1100 -3050 -1000 -2950
rect -850 -3000 -800 -2950
rect 1000 -2950 1100 -2850
rect 1950 -2450 2050 -2350
rect 1950 -2650 2050 -2550
rect 1950 -2850 2050 -2750
rect 1950 -3050 2050 -2950
rect -1100 -3250 -1000 -3150
rect 1950 -3250 2050 -3150
rect -17000 -14000 -9000 -6000
rect -4000 -14000 4000 -6000
rect 9000 -14000 17000 -6000
<< metal1 >>
rect -18000 12000 -8000 13000
rect -18000 4000 -17000 12000
rect -9000 4000 -8000 12000
rect -18000 3000 -8000 4000
rect -5000 12000 5000 13000
rect -5000 4000 -4000 12000
rect 4000 4000 5000 12000
rect -5000 3000 5000 4000
rect 8000 12000 18000 13000
rect 8000 4000 9000 12000
rect 17000 4000 18000 12000
rect 8000 3000 18000 4000
rect -15000 1000 -11000 3000
rect -100 1550 1800 3000
rect 12650 2450 14050 3000
rect 300 1500 1400 1550
rect 300 1350 800 1500
rect 950 1350 1400 1500
rect 300 1300 1400 1350
rect 12650 1250 12700 2450
rect 14000 1250 14050 2450
rect 12650 1200 14050 1250
rect -1150 1050 -950 1100
rect 1900 1050 2100 1100
rect -1150 1000 -1100 1050
rect -15000 950 -1100 1000
rect -1000 950 -950 1050
rect -15000 850 -950 950
rect -500 1000 -350 1050
rect -500 950 -450 1000
rect -400 950 -350 1000
rect -500 900 -350 950
rect 1900 950 1950 1050
rect 2050 1000 2100 1050
rect 2050 950 15000 1000
rect -15000 750 -1100 850
rect -1000 750 -950 850
rect -15000 650 -950 750
rect -900 800 -700 850
rect 500 800 700 850
rect 1100 800 1550 900
rect 1900 850 15000 950
rect 1900 800 1950 850
rect -900 700 -850 800
rect -750 700 -700 800
rect -900 650 -700 700
rect 50 700 550 800
rect 650 700 1200 800
rect 1450 750 1950 800
rect 2050 750 15000 850
rect 1450 700 15000 750
rect -15000 550 -1100 650
rect -1000 550 -950 650
rect -15000 450 -950 550
rect -800 600 -700 650
rect -150 600 0 650
rect 50 600 150 700
rect 500 650 700 700
rect 1250 650 1400 700
rect -800 550 -100 600
rect -50 550 150 600
rect 1250 600 1300 650
rect 1350 600 1400 650
rect 1250 550 1400 600
rect 1900 650 15000 700
rect 1900 550 1950 650
rect 2050 550 15000 650
rect -800 500 150 550
rect 1900 450 15000 550
rect -15000 350 -1100 450
rect -1000 350 -950 450
rect -15000 250 -950 350
rect -700 400 -500 450
rect 0 400 200 450
rect -700 300 -650 400
rect -550 300 50 400
rect 150 300 200 400
rect -700 250 -500 300
rect 0 250 200 300
rect 500 400 700 450
rect 1200 400 1400 450
rect 500 300 550 400
rect 650 300 1250 400
rect 1350 300 1400 400
rect 500 250 700 300
rect 1200 250 1400 300
rect 1900 350 1950 450
rect 2050 350 15000 450
rect 1900 250 15000 350
rect -15000 150 -1100 250
rect -1000 150 -950 250
rect 1900 150 1950 250
rect 2050 150 15000 250
rect -15000 50 -950 150
rect -15000 -50 -1100 50
rect -1000 -50 -950 50
rect -750 100 450 150
rect -750 50 -700 100
rect -650 50 350 100
rect 400 50 450 100
rect -750 0 -600 50
rect 300 0 450 50
rect 800 100 950 150
rect 800 50 850 100
rect 900 50 950 100
rect 800 0 950 50
rect 1550 100 1700 150
rect 1550 50 1600 100
rect 1650 50 1700 100
rect 1550 0 1700 50
rect 1900 50 15000 150
rect 1900 -50 1950 50
rect 2050 -50 15000 50
rect -15000 -150 -950 -50
rect -15000 -250 -1100 -150
rect -1000 -250 -950 -150
rect -900 -100 -700 -50
rect -900 -200 -850 -100
rect -750 -200 -700 -100
rect -900 -250 -700 -200
rect -450 -100 -250 -50
rect -450 -200 -400 -100
rect -300 -200 -250 -100
rect -450 -250 -250 -200
rect 0 -100 200 -50
rect 0 -200 50 -100
rect 150 -200 200 -100
rect 0 -250 200 -200
rect 500 -100 700 -50
rect 500 -200 550 -100
rect 650 -200 700 -100
rect 500 -250 700 -200
rect 950 -100 1150 -50
rect 1650 -100 1850 -50
rect 950 -200 1000 -100
rect 1100 -200 1150 -100
rect 950 -250 1150 -200
rect 1200 -150 1350 -100
rect 1200 -200 1250 -150
rect 1300 -200 1350 -150
rect 1200 -250 1350 -200
rect 1650 -200 1700 -100
rect 1800 -200 1850 -100
rect 1650 -250 1850 -200
rect 1900 -150 15000 -50
rect 1900 -250 1950 -150
rect 2050 -250 15000 -150
rect -15000 -350 -950 -250
rect -15000 -450 -1100 -350
rect -1000 -450 -950 -350
rect -15000 -550 -950 -450
rect -850 -550 -750 -250
rect -400 -550 -300 -250
rect 50 -550 150 -250
rect 550 -350 650 -250
rect 250 -450 650 -350
rect 550 -550 650 -450
rect -15000 -650 -1100 -550
rect -1000 -650 -950 -550
rect -15000 -750 -950 -650
rect -900 -600 -700 -550
rect -900 -700 -850 -600
rect -750 -700 -700 -600
rect -900 -750 -700 -700
rect -450 -600 -250 -550
rect -450 -700 -400 -600
rect -300 -700 -250 -600
rect -450 -750 -250 -700
rect 0 -600 200 -550
rect 500 -600 700 -550
rect 0 -700 50 -600
rect 150 -700 550 -600
rect 650 -700 700 -600
rect 0 -750 200 -700
rect 500 -750 700 -700
rect -15000 -850 -1100 -750
rect -1000 -850 -950 -750
rect -600 -850 -450 -800
rect -15000 -950 -950 -850
rect -15000 -1050 -1100 -950
rect -1000 -1050 -950 -950
rect -15000 -1150 -950 -1050
rect -15000 -1250 -1100 -1150
rect -1000 -1250 -950 -1150
rect -15000 -1350 -950 -1250
rect -15000 -1450 -1100 -1350
rect -1000 -1450 -950 -1350
rect -15000 -1550 -950 -1450
rect -15000 -1650 -1100 -1550
rect -1000 -1650 -950 -1550
rect -15000 -1750 -950 -1650
rect -15000 -1850 -1100 -1750
rect -1000 -1850 -950 -1750
rect -15000 -1950 -950 -1850
rect -15000 -2050 -1100 -1950
rect -1000 -2050 -950 -1950
rect -15000 -2150 -950 -2050
rect -15000 -2250 -1100 -2150
rect -1000 -2250 -950 -2150
rect -15000 -2350 -950 -2250
rect -15000 -2450 -1100 -2350
rect -1000 -2450 -950 -2350
rect -15000 -2550 -950 -2450
rect -15000 -2650 -1100 -2550
rect -1000 -2650 -950 -2550
rect -15000 -2750 -950 -2650
rect -15000 -2850 -1100 -2750
rect -1000 -2850 -950 -2750
rect -15000 -2950 -950 -2850
rect -15000 -3000 -1100 -2950
rect -1150 -3050 -1100 -3000
rect -1000 -3050 -950 -2950
rect -900 -900 -750 -850
rect -900 -950 -850 -900
rect -800 -950 -750 -900
rect -600 -900 -550 -850
rect -500 -900 -450 -850
rect -600 -950 -450 -900
rect 100 -850 250 -800
rect 1000 -850 1100 -250
rect 1900 -350 15000 -250
rect 1900 -450 1950 -350
rect 2050 -450 15000 -350
rect 1900 -550 15000 -450
rect 1250 -600 1400 -550
rect 1250 -650 1300 -600
rect 1350 -650 1400 -600
rect 1900 -650 1950 -550
rect 2050 -650 15000 -550
rect 1250 -700 1400 -650
rect 1450 -700 1600 -650
rect 100 -900 150 -850
rect 200 -900 1100 -850
rect 100 -950 1100 -900
rect 1450 -750 1500 -700
rect 1550 -750 1600 -700
rect 1450 -800 1600 -750
rect 1900 -750 15000 -650
rect -900 -1000 -750 -950
rect -900 -2450 -800 -1000
rect -700 -1250 -500 -1200
rect 700 -1250 900 -1200
rect -700 -1350 -650 -1250
rect -550 -1350 750 -1250
rect 850 -1350 900 -1250
rect 1450 -1350 1550 -800
rect 1650 -850 1800 -800
rect 1650 -900 1700 -850
rect 1750 -900 1800 -850
rect 1650 -950 1800 -900
rect 1900 -850 1950 -750
rect 2050 -850 15000 -750
rect 1900 -950 15000 -850
rect 1900 -1050 1950 -950
rect 2050 -1050 15000 -950
rect 1900 -1150 15000 -1050
rect 1900 -1250 1950 -1150
rect 2050 -1250 15000 -1150
rect -700 -1400 -500 -1350
rect 700 -1400 900 -1350
rect 1400 -1450 1550 -1350
rect 1650 -1350 1800 -1300
rect 1650 -1400 1700 -1350
rect 1750 -1400 1800 -1350
rect 1650 -1450 1800 -1400
rect 250 -1500 450 -1450
rect 250 -1600 300 -1500
rect 400 -1600 450 -1500
rect 250 -1650 450 -1600
rect 300 -2000 400 -1650
rect 1400 -2000 1500 -1450
rect 1700 -1700 1800 -1450
rect 1900 -1350 15000 -1250
rect 1900 -1450 1950 -1350
rect 2050 -1450 15000 -1350
rect 1900 -1550 15000 -1450
rect 1900 -1650 1950 -1550
rect 2050 -1650 15000 -1550
rect 1650 -1750 1850 -1700
rect 1650 -1850 1700 -1750
rect 1800 -1850 1850 -1750
rect 1650 -1900 1850 -1850
rect 1900 -1750 15000 -1650
rect 1900 -1850 1950 -1750
rect 2050 -1850 15000 -1750
rect -700 -2050 -550 -2000
rect -700 -2100 -650 -2050
rect -600 -2100 -550 -2050
rect -700 -2150 -550 -2100
rect -400 -2050 -250 -2000
rect -400 -2100 -350 -2050
rect -300 -2100 -250 -2050
rect -400 -2150 -250 -2100
rect -200 -2050 400 -2000
rect 700 -2050 850 -2000
rect -200 -2100 -150 -2050
rect -100 -2100 400 -2050
rect 450 -2100 750 -2050
rect 800 -2100 850 -2050
rect -200 -2150 -50 -2100
rect 450 -2150 850 -2100
rect 1350 -2050 1500 -2000
rect 1350 -2100 1400 -2050
rect 1450 -2100 1500 -2050
rect -400 -2450 -300 -2150
rect 50 -2250 250 -2200
rect 450 -2250 550 -2150
rect 50 -2350 100 -2250
rect 200 -2350 550 -2250
rect 50 -2400 250 -2350
rect -900 -2550 -300 -2450
rect 1350 -2500 1500 -2100
rect -900 -2900 -800 -2550
rect 0 -2700 1500 -2500
rect 1900 -1950 15000 -1850
rect 1900 -2050 1950 -1950
rect 2050 -2050 15000 -1950
rect 1900 -2150 15000 -2050
rect 1900 -2250 1950 -2150
rect 2050 -2250 15000 -2150
rect 1900 -2350 15000 -2250
rect 1900 -2450 1950 -2350
rect 2050 -2450 15000 -2350
rect 1900 -2550 15000 -2450
rect 1900 -2650 1950 -2550
rect 2050 -2650 15000 -2550
rect -900 -2950 -750 -2900
rect -900 -3000 -850 -2950
rect -800 -3000 -750 -2950
rect -900 -3050 -750 -3000
rect -1150 -3150 -950 -3050
rect -1150 -3250 -1100 -3150
rect -1000 -3250 -950 -3150
rect -1150 -3300 -950 -3250
rect 0 -3700 200 -2700
rect 1900 -2750 15000 -2650
rect 850 -2850 1250 -2800
rect 850 -2950 1000 -2850
rect 1100 -2950 1250 -2850
rect 850 -3350 1250 -2950
rect 1900 -2850 1950 -2750
rect 2050 -2850 15000 -2750
rect 1900 -2950 15000 -2850
rect 1900 -3050 1950 -2950
rect 2050 -3000 15000 -2950
rect 2050 -3050 2100 -3000
rect 1900 -3150 2100 -3050
rect 1900 -3250 1950 -3150
rect 2050 -3250 2100 -3150
rect 1900 -3300 2100 -3250
rect -10000 -4550 200 -3700
rect -10000 -5000 -9050 -4550
rect 650 -5000 1450 -3350
rect 11000 -5000 15000 -3000
rect -18000 -6000 -8000 -5000
rect -18000 -14000 -17000 -6000
rect -9000 -14000 -8000 -6000
rect -18000 -15000 -8000 -14000
rect -5000 -6000 5000 -5000
rect -5000 -14000 -4000 -6000
rect 4000 -14000 5000 -6000
rect -5000 -15000 5000 -14000
rect 8000 -6000 18000 -5000
rect 8000 -14000 9000 -6000
rect 17000 -14000 18000 -6000
rect 8000 -15000 18000 -14000
<< via1 >>
rect 800 1350 950 1500
rect 12700 1250 14000 2450
rect -450 950 -400 1000
rect 1300 600 1350 650
rect -700 50 -650 100
rect 850 50 900 100
rect 1600 50 1650 100
rect 550 -200 650 -100
rect 1250 -200 1300 -150
rect -850 -700 -750 -600
rect 50 -700 150 -600
rect -550 -900 -500 -850
rect 1300 -650 1350 -600
rect 1500 -750 1550 -700
rect 750 -1350 850 -1250
rect 1700 -900 1750 -850
rect 1950 -1250 2050 -1150
rect -650 -2100 -600 -2050
<< metal2 >>
rect 3500 2450 14050 2500
rect 3500 2000 12700 2450
rect 750 1500 1000 1550
rect 750 1350 800 1500
rect 950 1350 1000 1500
rect 2200 1350 12700 2000
rect 750 1300 1000 1350
rect 1750 1250 12700 1350
rect 14000 1250 14050 2450
rect 1750 1200 14050 1250
rect -500 1000 -350 1050
rect -500 950 -450 1000
rect -400 950 1550 1000
rect -500 900 1550 950
rect 1250 650 1400 700
rect 1250 600 1300 650
rect 1350 600 1400 650
rect 1250 550 1400 600
rect -750 100 -600 150
rect -750 50 -700 100
rect -650 50 -600 100
rect -750 0 -600 50
rect 800 100 950 150
rect 800 50 850 100
rect 900 50 950 100
rect 1250 50 1350 550
rect 1450 300 1550 900
rect 800 0 950 50
rect 1000 -50 1350 50
rect 1400 200 1550 300
rect 1400 -50 1500 200
rect 1750 150 1900 1200
rect 1550 100 1900 150
rect 1550 50 1600 100
rect 1650 50 1900 100
rect 1550 0 1900 50
rect 500 -100 700 -50
rect 500 -200 550 -100
rect 650 -200 700 -100
rect 500 -250 700 -200
rect 900 -150 1100 -50
rect 1200 -150 1350 -100
rect 1400 -150 1550 -50
rect 900 -550 1000 -150
rect 1200 -200 1250 -150
rect 1300 -200 1350 -150
rect 1200 -250 1350 -200
rect -900 -600 -700 -550
rect 0 -600 200 -550
rect -900 -700 -850 -600
rect -750 -700 50 -600
rect 150 -700 200 -600
rect 900 -600 1400 -550
rect 900 -650 1300 -600
rect 1350 -650 1400 -600
rect 1250 -700 1400 -650
rect 1450 -650 1550 -150
rect 1450 -700 1600 -650
rect -900 -750 -700 -700
rect 0 -750 200 -700
rect 1450 -750 1500 -700
rect 1550 -750 1600 -700
rect 1450 -800 1600 -750
rect -600 -850 -450 -800
rect 1650 -850 1800 -800
rect -600 -900 -550 -850
rect -500 -900 1700 -850
rect 1750 -900 1800 -850
rect -600 -950 1800 -900
rect 1900 -1150 2100 -1100
rect 1900 -1200 1950 -1150
rect 700 -1250 1950 -1200
rect 2050 -1250 2100 -1150
rect 700 -1350 750 -1250
rect 850 -1300 2100 -1250
rect 850 -1350 900 -1300
rect 700 -1400 900 -1350
rect -700 -2050 -550 -2000
rect -700 -2100 -650 -2050
rect -600 -2100 -550 -2050
rect -700 -2150 -550 -2100
<< via2 >>
rect 800 1350 950 1500
rect -700 50 -650 100
rect 850 50 900 100
rect 550 -200 650 -100
rect 1250 -200 1300 -150
rect -650 -2100 -600 -2050
<< metal3 >>
rect 750 1500 1000 1550
rect 750 1350 800 1500
rect 950 1350 1000 1500
rect 750 1300 1000 1350
rect -750 100 -600 150
rect -750 50 -700 100
rect -650 50 -600 100
rect -750 0 -600 50
rect 800 100 950 1300
rect 800 50 850 100
rect 900 50 950 100
rect 800 0 950 50
rect -700 -2000 -600 0
rect 500 -100 700 -50
rect 1250 -100 1350 -50
rect 500 -200 550 -100
rect 650 -150 700 -100
rect 1200 -150 1350 -100
rect 650 -200 1250 -150
rect 1300 -200 1350 -150
rect 500 -250 1350 -200
rect -700 -2050 -550 -2000
rect -700 -2100 -650 -2050
rect -600 -2100 -550 -2050
rect -700 -2150 -550 -2100
<< labels >>
rlabel metal1 -18000 3000 -8000 13000 1 gnd
rlabel metal1 8000 -15000 18000 -5000 1 vdd
rlabel metal1 -5000 -15000 5000 -5000 1 out
rlabel metal1 -18000 -15000 -8000 -5000 1 clk
rlabel metal1 -5000 3000 5000 13000 1 inn
rlabel metal1 8000 3000 18000 13000 1 inp
rlabel locali -150 700 -50 800 1 net1
rlabel metal3 -750 0 -600 150 1 outn
rlabel locali -400 -50 -300 50 1 outp
rlabel locali 1000 50 1100 150 1 net3
rlabel locali 1700 -400 1800 -300 1 net2
rlabel locali 1050 550 1150 650 1 clkb
rlabel locali 750 -450 850 -350 1 net4
rlabel locali -400 -1600 -300 -1500 1 net5
rlabel locali 100 -2150 200 -2050 1 net7
rlabel metal1 -400 -2150 -250 -2000 1 net6
rlabel locali -200 -2550 -100 -2450 1 net8
<< end >>
